module hazard_unit(

)

endmodule