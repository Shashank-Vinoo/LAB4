module control_hazard_unit(

)

endmodule