module data_hazard_unit (

)

endmodule